* File: total.pex.spi
* Created: Thu Dec 28 19:20:33 2023
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "total.pex.spi.pex"
.subckt total  F_4_INV F_4 F_2 F_2_INV F_32_INV F_32 F_16 F_16_INV F_8 F_8_INV
+ F_64 F_64_INV EN CLK_IN RST GND VDD WL<5> WL<1> WL<7> WL<3> WL<4> WL<0> WL<6>
+ WL<2> BL<5> BL<1> BL<7> BL<3> BL<4> BL<0> BL<6> BL<2>
* 
* BL<2>	BL<2>
* BL<6>	BL<6>
* BL<0>	BL<0>
* BL<4>	BL<4>
* BL<3>	BL<3>
* BL<7>	BL<7>
* BL<1>	BL<1>
* BL<5>	BL<5>
* WL<2>	WL<2>
* WL<6>	WL<6>
* WL<0>	WL<0>
* WL<4>	WL<4>
* WL<3>	WL<3>
* WL<7>	WL<7>
* WL<1>	WL<1>
* WL<5>	WL<5>
* VDD	VDD
* GND	GND
* RST	RST
* CLK_IN	CLK_IN
* EN	EN
* F_64_INV	F_64_INV
* F_64	F_64
* F_8_INV	F_8_INV
* F_8	F_8
* F_16_INV	F_16_INV
* F_16	F_16
* F_32	F_32
* F_32_INV	F_32_INV
* F_2_INV	F_2_INV
* F_2	F_2
* F_4	F_4
* F_4_INV	F_4_INV
mXI2.XI5.MMN1 N_XI2.XI5.NET27_XI2.XI5.MMN1_d N_F_64_XI2.XI5.MMN1_g
+ N_GND_XI2.XI5.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI5.MMN2 N_XI2.XI5.NET28_XI2.XI5.MMN2_d N_F_32_INV_XI2.XI5.MMN2_g
+ N_XI2.XI5.NET27_XI2.XI5.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI5.MMN3 N_XI2.XI5.NET16_XI2.XI5.MMN3_d N_F_16_XI2.XI5.MMN3_g
+ N_XI2.XI5.NET28_XI2.XI5.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI5.MMinv2 N_WL<5>_XI2.XI5.MMinv2_d N_XI2.XI5.NET16_XI2.XI5.MMinv2_g
+ N_GND_XI2.XI5.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI5.MMinv2@4 N_WL<5>_XI2.XI5.MMinv2@4_d N_XI2.XI5.NET16_XI2.XI5.MMinv2@4_g
+ N_GND_XI2.XI5.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMinv2@3 N_WL<5>_XI2.XI5.MMinv2@3_d N_XI2.XI5.NET16_XI2.XI5.MMinv2@3_g
+ N_GND_XI2.XI5.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMinv2@2 N_WL<5>_XI2.XI5.MMinv2@2_d N_XI2.XI5.NET16_XI2.XI5.MMinv2@2_g
+ N_GND_XI2.XI5.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI5.MMP1 N_XI2.XI5.NET16_XI2.XI5.MMP1_d N_F_64_XI2.XI5.MMP1_g
+ N_VDD_XI2.XI5.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI5.MMP2 N_XI2.XI5.NET16_XI2.XI5.MMP2_d N_F_32_INV_XI2.XI5.MMP2_g
+ N_VDD_XI2.XI5.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMP3 N_XI2.XI5.NET16_XI2.XI5.MMP3_d N_F_16_XI2.XI5.MMP3_g
+ N_VDD_XI2.XI5.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI5.MMen N_XI2.XI5.NET16_XI2.XI5.MMen_d N_EN_XI2.XI5.MMen_g
+ N_VDD_XI2.XI5.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI5.MMinv1 N_WL<5>_XI2.XI5.MMinv1_d N_XI2.XI5.NET16_XI2.XI5.MMinv1_g
+ N_VDD_XI2.XI5.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMinv1@4 N_WL<5>_XI2.XI5.MMinv1@4_d N_XI2.XI5.NET16_XI2.XI5.MMinv1@4_g
+ N_VDD_XI2.XI5.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMinv1@3 N_WL<5>_XI2.XI5.MMinv1@3_d N_XI2.XI5.NET16_XI2.XI5.MMinv1@3_g
+ N_VDD_XI2.XI5.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI5.MMinv1@2 N_WL<5>_XI2.XI5.MMinv1@2_d N_XI2.XI5.NET16_XI2.XI5.MMinv1@2_g
+ N_VDD_XI2.XI5.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI1.MMN1 N_XI2.XI1.NET27_XI2.XI1.MMN1_d N_F_64_INV_XI2.XI1.MMN1_g
+ N_GND_XI2.XI1.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI1.MMN2 N_XI2.XI1.NET28_XI2.XI1.MMN2_d N_F_32_INV_XI2.XI1.MMN2_g
+ N_XI2.XI1.NET27_XI2.XI1.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI1.MMN3 N_XI2.XI1.NET16_XI2.XI1.MMN3_d N_F_16_XI2.XI1.MMN3_g
+ N_XI2.XI1.NET28_XI2.XI1.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI1.MMinv2 N_WL<1>_XI2.XI1.MMinv2_d N_XI2.XI1.NET16_XI2.XI1.MMinv2_g
+ N_GND_XI2.XI1.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI1.MMinv2@4 N_WL<1>_XI2.XI1.MMinv2@4_d N_XI2.XI1.NET16_XI2.XI1.MMinv2@4_g
+ N_GND_XI2.XI1.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMinv2@3 N_WL<1>_XI2.XI1.MMinv2@3_d N_XI2.XI1.NET16_XI2.XI1.MMinv2@3_g
+ N_GND_XI2.XI1.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMinv2@2 N_WL<1>_XI2.XI1.MMinv2@2_d N_XI2.XI1.NET16_XI2.XI1.MMinv2@2_g
+ N_GND_XI2.XI1.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI1.MMP1 N_XI2.XI1.NET16_XI2.XI1.MMP1_d N_F_64_INV_XI2.XI1.MMP1_g
+ N_VDD_XI2.XI1.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI1.MMP2 N_XI2.XI1.NET16_XI2.XI1.MMP2_d N_F_32_INV_XI2.XI1.MMP2_g
+ N_VDD_XI2.XI1.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMP3 N_XI2.XI1.NET16_XI2.XI1.MMP3_d N_F_16_XI2.XI1.MMP3_g
+ N_VDD_XI2.XI1.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI1.MMen N_XI2.XI1.NET16_XI2.XI1.MMen_d N_EN_XI2.XI1.MMen_g
+ N_VDD_XI2.XI1.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI1.MMinv1 N_WL<1>_XI2.XI1.MMinv1_d N_XI2.XI1.NET16_XI2.XI1.MMinv1_g
+ N_VDD_XI2.XI1.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMinv1@4 N_WL<1>_XI2.XI1.MMinv1@4_d N_XI2.XI1.NET16_XI2.XI1.MMinv1@4_g
+ N_VDD_XI2.XI1.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMinv1@3 N_WL<1>_XI2.XI1.MMinv1@3_d N_XI2.XI1.NET16_XI2.XI1.MMinv1@3_g
+ N_VDD_XI2.XI1.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI1.MMinv1@2 N_WL<1>_XI2.XI1.MMinv1@2_d N_XI2.XI1.NET16_XI2.XI1.MMinv1@2_g
+ N_VDD_XI2.XI1.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI7.MMN1 N_XI2.XI7.NET27_XI2.XI7.MMN1_d N_F_64_XI2.XI7.MMN1_g
+ N_GND_XI2.XI7.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI7.MMN2 N_XI2.XI7.NET28_XI2.XI7.MMN2_d N_F_32_XI2.XI7.MMN2_g
+ N_XI2.XI7.NET27_XI2.XI7.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI7.MMN3 N_XI2.XI7.NET16_XI2.XI7.MMN3_d N_F_16_XI2.XI7.MMN3_g
+ N_XI2.XI7.NET28_XI2.XI7.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI7.MMinv2 N_WL<7>_XI2.XI7.MMinv2_d N_XI2.XI7.NET16_XI2.XI7.MMinv2_g
+ N_GND_XI2.XI7.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI7.MMinv2@4 N_WL<7>_XI2.XI7.MMinv2@4_d N_XI2.XI7.NET16_XI2.XI7.MMinv2@4_g
+ N_GND_XI2.XI7.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMinv2@3 N_WL<7>_XI2.XI7.MMinv2@3_d N_XI2.XI7.NET16_XI2.XI7.MMinv2@3_g
+ N_GND_XI2.XI7.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMinv2@2 N_WL<7>_XI2.XI7.MMinv2@2_d N_XI2.XI7.NET16_XI2.XI7.MMinv2@2_g
+ N_GND_XI2.XI7.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI7.MMP1 N_XI2.XI7.NET16_XI2.XI7.MMP1_d N_F_64_XI2.XI7.MMP1_g
+ N_VDD_XI2.XI7.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI7.MMP2 N_XI2.XI7.NET16_XI2.XI7.MMP2_d N_F_32_XI2.XI7.MMP2_g
+ N_VDD_XI2.XI7.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMP3 N_XI2.XI7.NET16_XI2.XI7.MMP3_d N_F_16_XI2.XI7.MMP3_g
+ N_VDD_XI2.XI7.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI7.MMen N_XI2.XI7.NET16_XI2.XI7.MMen_d N_EN_XI2.XI7.MMen_g
+ N_VDD_XI2.XI7.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI7.MMinv1 N_WL<7>_XI2.XI7.MMinv1_d N_XI2.XI7.NET16_XI2.XI7.MMinv1_g
+ N_VDD_XI2.XI7.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMinv1@4 N_WL<7>_XI2.XI7.MMinv1@4_d N_XI2.XI7.NET16_XI2.XI7.MMinv1@4_g
+ N_VDD_XI2.XI7.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMinv1@3 N_WL<7>_XI2.XI7.MMinv1@3_d N_XI2.XI7.NET16_XI2.XI7.MMinv1@3_g
+ N_VDD_XI2.XI7.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI7.MMinv1@2 N_WL<7>_XI2.XI7.MMinv1@2_d N_XI2.XI7.NET16_XI2.XI7.MMinv1@2_g
+ N_VDD_XI2.XI7.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI3.MMN1 N_XI2.XI3.NET27_XI2.XI3.MMN1_d N_F_64_INV_XI2.XI3.MMN1_g
+ N_GND_XI2.XI3.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI3.MMN2 N_XI2.XI3.NET28_XI2.XI3.MMN2_d N_F_32_XI2.XI3.MMN2_g
+ N_XI2.XI3.NET27_XI2.XI3.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI3.MMN3 N_XI2.XI3.NET16_XI2.XI3.MMN3_d N_F_16_XI2.XI3.MMN3_g
+ N_XI2.XI3.NET28_XI2.XI3.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI3.MMinv2 N_WL<3>_XI2.XI3.MMinv2_d N_XI2.XI3.NET16_XI2.XI3.MMinv2_g
+ N_GND_XI2.XI3.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI3.MMinv2@4 N_WL<3>_XI2.XI3.MMinv2@4_d N_XI2.XI3.NET16_XI2.XI3.MMinv2@4_g
+ N_GND_XI2.XI3.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMinv2@3 N_WL<3>_XI2.XI3.MMinv2@3_d N_XI2.XI3.NET16_XI2.XI3.MMinv2@3_g
+ N_GND_XI2.XI3.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMinv2@2 N_WL<3>_XI2.XI3.MMinv2@2_d N_XI2.XI3.NET16_XI2.XI3.MMinv2@2_g
+ N_GND_XI2.XI3.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI3.MMP1 N_XI2.XI3.NET16_XI2.XI3.MMP1_d N_F_64_INV_XI2.XI3.MMP1_g
+ N_VDD_XI2.XI3.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI3.MMP2 N_XI2.XI3.NET16_XI2.XI3.MMP2_d N_F_32_XI2.XI3.MMP2_g
+ N_VDD_XI2.XI3.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMP3 N_XI2.XI3.NET16_XI2.XI3.MMP3_d N_F_16_XI2.XI3.MMP3_g
+ N_VDD_XI2.XI3.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI3.MMen N_XI2.XI3.NET16_XI2.XI3.MMen_d N_EN_XI2.XI3.MMen_g
+ N_VDD_XI2.XI3.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI3.MMinv1 N_WL<3>_XI2.XI3.MMinv1_d N_XI2.XI3.NET16_XI2.XI3.MMinv1_g
+ N_VDD_XI2.XI3.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMinv1@4 N_WL<3>_XI2.XI3.MMinv1@4_d N_XI2.XI3.NET16_XI2.XI3.MMinv1@4_g
+ N_VDD_XI2.XI3.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMinv1@3 N_WL<3>_XI2.XI3.MMinv1@3_d N_XI2.XI3.NET16_XI2.XI3.MMinv1@3_g
+ N_VDD_XI2.XI3.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI3.MMinv1@2 N_WL<3>_XI2.XI3.MMinv1@2_d N_XI2.XI3.NET16_XI2.XI3.MMinv1@2_g
+ N_VDD_XI2.XI3.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI4.MMN1 N_XI2.XI4.NET27_XI2.XI4.MMN1_d N_F_64_XI2.XI4.MMN1_g
+ N_GND_XI2.XI4.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI4.MMN2 N_XI2.XI4.NET28_XI2.XI4.MMN2_d N_F_32_INV_XI2.XI4.MMN2_g
+ N_XI2.XI4.NET27_XI2.XI4.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI4.MMN3 N_XI2.XI4.NET16_XI2.XI4.MMN3_d N_F_16_INV_XI2.XI4.MMN3_g
+ N_XI2.XI4.NET28_XI2.XI4.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI4.MMinv2 N_WL<4>_XI2.XI4.MMinv2_d N_XI2.XI4.NET16_XI2.XI4.MMinv2_g
+ N_GND_XI2.XI4.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI4.MMinv2@4 N_WL<4>_XI2.XI4.MMinv2@4_d N_XI2.XI4.NET16_XI2.XI4.MMinv2@4_g
+ N_GND_XI2.XI4.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMinv2@3 N_WL<4>_XI2.XI4.MMinv2@3_d N_XI2.XI4.NET16_XI2.XI4.MMinv2@3_g
+ N_GND_XI2.XI4.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMinv2@2 N_WL<4>_XI2.XI4.MMinv2@2_d N_XI2.XI4.NET16_XI2.XI4.MMinv2@2_g
+ N_GND_XI2.XI4.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI4.MMP1 N_XI2.XI4.NET16_XI2.XI4.MMP1_d N_F_64_XI2.XI4.MMP1_g
+ N_VDD_XI2.XI4.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI4.MMP2 N_XI2.XI4.NET16_XI2.XI4.MMP2_d N_F_32_INV_XI2.XI4.MMP2_g
+ N_VDD_XI2.XI4.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMP3 N_XI2.XI4.NET16_XI2.XI4.MMP3_d N_F_16_INV_XI2.XI4.MMP3_g
+ N_VDD_XI2.XI4.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI4.MMen N_XI2.XI4.NET16_XI2.XI4.MMen_d N_EN_XI2.XI4.MMen_g
+ N_VDD_XI2.XI4.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI4.MMinv1 N_WL<4>_XI2.XI4.MMinv1_d N_XI2.XI4.NET16_XI2.XI4.MMinv1_g
+ N_VDD_XI2.XI4.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMinv1@4 N_WL<4>_XI2.XI4.MMinv1@4_d N_XI2.XI4.NET16_XI2.XI4.MMinv1@4_g
+ N_VDD_XI2.XI4.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMinv1@3 N_WL<4>_XI2.XI4.MMinv1@3_d N_XI2.XI4.NET16_XI2.XI4.MMinv1@3_g
+ N_VDD_XI2.XI4.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI4.MMinv1@2 N_WL<4>_XI2.XI4.MMinv1@2_d N_XI2.XI4.NET16_XI2.XI4.MMinv1@2_g
+ N_VDD_XI2.XI4.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI0.MMN1 N_XI2.XI0.NET27_XI2.XI0.MMN1_d N_F_64_INV_XI2.XI0.MMN1_g
+ N_GND_XI2.XI0.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI0.MMN2 N_XI2.XI0.NET28_XI2.XI0.MMN2_d N_F_32_INV_XI2.XI0.MMN2_g
+ N_XI2.XI0.NET27_XI2.XI0.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI0.MMN3 N_XI2.XI0.NET16_XI2.XI0.MMN3_d N_F_16_INV_XI2.XI0.MMN3_g
+ N_XI2.XI0.NET28_XI2.XI0.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI0.MMinv2 N_WL<0>_XI2.XI0.MMinv2_d N_XI2.XI0.NET16_XI2.XI0.MMinv2_g
+ N_GND_XI2.XI0.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI0.MMinv2@4 N_WL<0>_XI2.XI0.MMinv2@4_d N_XI2.XI0.NET16_XI2.XI0.MMinv2@4_g
+ N_GND_XI2.XI0.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMinv2@3 N_WL<0>_XI2.XI0.MMinv2@3_d N_XI2.XI0.NET16_XI2.XI0.MMinv2@3_g
+ N_GND_XI2.XI0.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMinv2@2 N_WL<0>_XI2.XI0.MMinv2@2_d N_XI2.XI0.NET16_XI2.XI0.MMinv2@2_g
+ N_GND_XI2.XI0.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI0.MMP1 N_XI2.XI0.NET16_XI2.XI0.MMP1_d N_F_64_INV_XI2.XI0.MMP1_g
+ N_VDD_XI2.XI0.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI0.MMP2 N_XI2.XI0.NET16_XI2.XI0.MMP2_d N_F_32_INV_XI2.XI0.MMP2_g
+ N_VDD_XI2.XI0.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMP3 N_XI2.XI0.NET16_XI2.XI0.MMP3_d N_F_16_INV_XI2.XI0.MMP3_g
+ N_VDD_XI2.XI0.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI0.MMen N_XI2.XI0.NET16_XI2.XI0.MMen_d N_EN_XI2.XI0.MMen_g
+ N_VDD_XI2.XI0.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI0.MMinv1 N_WL<0>_XI2.XI0.MMinv1_d N_XI2.XI0.NET16_XI2.XI0.MMinv1_g
+ N_VDD_XI2.XI0.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMinv1@4 N_WL<0>_XI2.XI0.MMinv1@4_d N_XI2.XI0.NET16_XI2.XI0.MMinv1@4_g
+ N_VDD_XI2.XI0.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMinv1@3 N_WL<0>_XI2.XI0.MMinv1@3_d N_XI2.XI0.NET16_XI2.XI0.MMinv1@3_g
+ N_VDD_XI2.XI0.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI0.MMinv1@2 N_WL<0>_XI2.XI0.MMinv1@2_d N_XI2.XI0.NET16_XI2.XI0.MMinv1@2_g
+ N_VDD_XI2.XI0.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI6.MMN1 N_XI2.XI6.NET27_XI2.XI6.MMN1_d N_F_64_XI2.XI6.MMN1_g
+ N_GND_XI2.XI6.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI6.MMN2 N_XI2.XI6.NET28_XI2.XI6.MMN2_d N_F_32_XI2.XI6.MMN2_g
+ N_XI2.XI6.NET27_XI2.XI6.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI6.MMN3 N_XI2.XI6.NET16_XI2.XI6.MMN3_d N_F_16_INV_XI2.XI6.MMN3_g
+ N_XI2.XI6.NET28_XI2.XI6.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI6.MMinv2 N_WL<6>_XI2.XI6.MMinv2_d N_XI2.XI6.NET16_XI2.XI6.MMinv2_g
+ N_GND_XI2.XI6.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI6.MMinv2@4 N_WL<6>_XI2.XI6.MMinv2@4_d N_XI2.XI6.NET16_XI2.XI6.MMinv2@4_g
+ N_GND_XI2.XI6.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMinv2@3 N_WL<6>_XI2.XI6.MMinv2@3_d N_XI2.XI6.NET16_XI2.XI6.MMinv2@3_g
+ N_GND_XI2.XI6.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMinv2@2 N_WL<6>_XI2.XI6.MMinv2@2_d N_XI2.XI6.NET16_XI2.XI6.MMinv2@2_g
+ N_GND_XI2.XI6.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI6.MMP1 N_XI2.XI6.NET16_XI2.XI6.MMP1_d N_F_64_XI2.XI6.MMP1_g
+ N_VDD_XI2.XI6.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI6.MMP2 N_XI2.XI6.NET16_XI2.XI6.MMP2_d N_F_32_XI2.XI6.MMP2_g
+ N_VDD_XI2.XI6.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMP3 N_XI2.XI6.NET16_XI2.XI6.MMP3_d N_F_16_INV_XI2.XI6.MMP3_g
+ N_VDD_XI2.XI6.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI6.MMen N_XI2.XI6.NET16_XI2.XI6.MMen_d N_EN_XI2.XI6.MMen_g
+ N_VDD_XI2.XI6.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI6.MMinv1 N_WL<6>_XI2.XI6.MMinv1_d N_XI2.XI6.NET16_XI2.XI6.MMinv1_g
+ N_VDD_XI2.XI6.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMinv1@4 N_WL<6>_XI2.XI6.MMinv1@4_d N_XI2.XI6.NET16_XI2.XI6.MMinv1@4_g
+ N_VDD_XI2.XI6.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMinv1@3 N_WL<6>_XI2.XI6.MMinv1@3_d N_XI2.XI6.NET16_XI2.XI6.MMinv1@3_g
+ N_VDD_XI2.XI6.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI6.MMinv1@2 N_WL<6>_XI2.XI6.MMinv1@2_d N_XI2.XI6.NET16_XI2.XI6.MMinv1@2_g
+ N_VDD_XI2.XI6.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI2.XI2.MMN1 N_XI2.XI2.NET27_XI2.XI2.MMN1_d N_F_64_INV_XI2.XI2.MMN1_g
+ N_GND_XI2.XI2.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI2.XI2.MMN2 N_XI2.XI2.NET28_XI2.XI2.MMN2_d N_F_32_XI2.XI2.MMN2_g
+ N_XI2.XI2.NET27_XI2.XI2.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI2.XI2.MMN3 N_XI2.XI2.NET16_XI2.XI2.MMN3_d N_F_16_INV_XI2.XI2.MMN3_g
+ N_XI2.XI2.NET28_XI2.XI2.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI2.XI2.MMinv2 N_WL<2>_XI2.XI2.MMinv2_d N_XI2.XI2.NET16_XI2.XI2.MMinv2_g
+ N_GND_XI2.XI2.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI2.MMinv2@4 N_WL<2>_XI2.XI2.MMinv2@4_d N_XI2.XI2.NET16_XI2.XI2.MMinv2@4_g
+ N_GND_XI2.XI2.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMinv2@3 N_WL<2>_XI2.XI2.MMinv2@3_d N_XI2.XI2.NET16_XI2.XI2.MMinv2@3_g
+ N_GND_XI2.XI2.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMinv2@2 N_WL<2>_XI2.XI2.MMinv2@2_d N_XI2.XI2.NET16_XI2.XI2.MMinv2@2_g
+ N_GND_XI2.XI2.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI2.XI2.MMP1 N_XI2.XI2.NET16_XI2.XI2.MMP1_d N_F_64_INV_XI2.XI2.MMP1_g
+ N_VDD_XI2.XI2.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI2.XI2.MMP2 N_XI2.XI2.NET16_XI2.XI2.MMP2_d N_F_32_XI2.XI2.MMP2_g
+ N_VDD_XI2.XI2.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMP3 N_XI2.XI2.NET16_XI2.XI2.MMP3_d N_F_16_INV_XI2.XI2.MMP3_g
+ N_VDD_XI2.XI2.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI2.XI2.MMen N_XI2.XI2.NET16_XI2.XI2.MMen_d N_EN_XI2.XI2.MMen_g
+ N_VDD_XI2.XI2.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI2.XI2.MMinv1 N_WL<2>_XI2.XI2.MMinv1_d N_XI2.XI2.NET16_XI2.XI2.MMinv1_g
+ N_VDD_XI2.XI2.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMinv1@4 N_WL<2>_XI2.XI2.MMinv1@4_d N_XI2.XI2.NET16_XI2.XI2.MMinv1@4_g
+ N_VDD_XI2.XI2.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMinv1@3 N_WL<2>_XI2.XI2.MMinv1@3_d N_XI2.XI2.NET16_XI2.XI2.MMinv1@3_g
+ N_VDD_XI2.XI2.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI2.XI2.MMinv1@2 N_WL<2>_XI2.XI2.MMinv1@2_d N_XI2.XI2.NET16_XI2.XI2.MMinv1@2_g
+ N_VDD_XI2.XI2.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI5.MMN1 N_XI1.XI5.NET27_XI1.XI5.MMN1_d N_F_8_XI1.XI5.MMN1_g
+ N_GND_XI1.XI5.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI5.MMN2 N_XI1.XI5.NET28_XI1.XI5.MMN2_d N_F_4_INV_XI1.XI5.MMN2_g
+ N_XI1.XI5.NET27_XI1.XI5.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI5.MMN3 N_XI1.XI5.NET16_XI1.XI5.MMN3_d N_F_2_XI1.XI5.MMN3_g
+ N_XI1.XI5.NET28_XI1.XI5.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI5.MMinv2 N_BL<5>_XI1.XI5.MMinv2_d N_XI1.XI5.NET16_XI1.XI5.MMinv2_g
+ N_GND_XI1.XI5.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI5.MMinv2@4 N_BL<5>_XI1.XI5.MMinv2@4_d N_XI1.XI5.NET16_XI1.XI5.MMinv2@4_g
+ N_GND_XI1.XI5.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMinv2@3 N_BL<5>_XI1.XI5.MMinv2@3_d N_XI1.XI5.NET16_XI1.XI5.MMinv2@3_g
+ N_GND_XI1.XI5.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMinv2@2 N_BL<5>_XI1.XI5.MMinv2@2_d N_XI1.XI5.NET16_XI1.XI5.MMinv2@2_g
+ N_GND_XI1.XI5.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI5.MMP1 N_XI1.XI5.NET16_XI1.XI5.MMP1_d N_F_8_XI1.XI5.MMP1_g
+ N_VDD_XI1.XI5.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI5.MMP2 N_XI1.XI5.NET16_XI1.XI5.MMP2_d N_F_4_INV_XI1.XI5.MMP2_g
+ N_VDD_XI1.XI5.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMP3 N_XI1.XI5.NET16_XI1.XI5.MMP3_d N_F_2_XI1.XI5.MMP3_g
+ N_VDD_XI1.XI5.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI5.MMen N_XI1.XI5.NET16_XI1.XI5.MMen_d N_EN_XI1.XI5.MMen_g
+ N_VDD_XI1.XI5.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI5.MMinv1 N_BL<5>_XI1.XI5.MMinv1_d N_XI1.XI5.NET16_XI1.XI5.MMinv1_g
+ N_VDD_XI1.XI5.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMinv1@4 N_BL<5>_XI1.XI5.MMinv1@4_d N_XI1.XI5.NET16_XI1.XI5.MMinv1@4_g
+ N_VDD_XI1.XI5.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMinv1@3 N_BL<5>_XI1.XI5.MMinv1@3_d N_XI1.XI5.NET16_XI1.XI5.MMinv1@3_g
+ N_VDD_XI1.XI5.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI5.MMinv1@2 N_BL<5>_XI1.XI5.MMinv1@2_d N_XI1.XI5.NET16_XI1.XI5.MMinv1@2_g
+ N_VDD_XI1.XI5.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI1.MMN1 N_XI1.XI1.NET27_XI1.XI1.MMN1_d N_F_8_INV_XI1.XI1.MMN1_g
+ N_GND_XI1.XI1.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI1.MMN2 N_XI1.XI1.NET28_XI1.XI1.MMN2_d N_F_4_INV_XI1.XI1.MMN2_g
+ N_XI1.XI1.NET27_XI1.XI1.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI1.MMN3 N_XI1.XI1.NET16_XI1.XI1.MMN3_d N_F_2_XI1.XI1.MMN3_g
+ N_XI1.XI1.NET28_XI1.XI1.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI1.MMinv2 N_BL<1>_XI1.XI1.MMinv2_d N_XI1.XI1.NET16_XI1.XI1.MMinv2_g
+ N_GND_XI1.XI1.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI1.MMinv2@4 N_BL<1>_XI1.XI1.MMinv2@4_d N_XI1.XI1.NET16_XI1.XI1.MMinv2@4_g
+ N_GND_XI1.XI1.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMinv2@3 N_BL<1>_XI1.XI1.MMinv2@3_d N_XI1.XI1.NET16_XI1.XI1.MMinv2@3_g
+ N_GND_XI1.XI1.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMinv2@2 N_BL<1>_XI1.XI1.MMinv2@2_d N_XI1.XI1.NET16_XI1.XI1.MMinv2@2_g
+ N_GND_XI1.XI1.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI1.MMP1 N_XI1.XI1.NET16_XI1.XI1.MMP1_d N_F_8_INV_XI1.XI1.MMP1_g
+ N_VDD_XI1.XI1.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI1.MMP2 N_XI1.XI1.NET16_XI1.XI1.MMP2_d N_F_4_INV_XI1.XI1.MMP2_g
+ N_VDD_XI1.XI1.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMP3 N_XI1.XI1.NET16_XI1.XI1.MMP3_d N_F_2_XI1.XI1.MMP3_g
+ N_VDD_XI1.XI1.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI1.MMen N_XI1.XI1.NET16_XI1.XI1.MMen_d N_EN_XI1.XI1.MMen_g
+ N_VDD_XI1.XI1.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI1.MMinv1 N_BL<1>_XI1.XI1.MMinv1_d N_XI1.XI1.NET16_XI1.XI1.MMinv1_g
+ N_VDD_XI1.XI1.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMinv1@4 N_BL<1>_XI1.XI1.MMinv1@4_d N_XI1.XI1.NET16_XI1.XI1.MMinv1@4_g
+ N_VDD_XI1.XI1.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMinv1@3 N_BL<1>_XI1.XI1.MMinv1@3_d N_XI1.XI1.NET16_XI1.XI1.MMinv1@3_g
+ N_VDD_XI1.XI1.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI1.MMinv1@2 N_BL<1>_XI1.XI1.MMinv1@2_d N_XI1.XI1.NET16_XI1.XI1.MMinv1@2_g
+ N_VDD_XI1.XI1.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI7.MMN1 N_XI1.XI7.NET27_XI1.XI7.MMN1_d N_F_8_XI1.XI7.MMN1_g
+ N_GND_XI1.XI7.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI7.MMN2 N_XI1.XI7.NET28_XI1.XI7.MMN2_d N_F_4_XI1.XI7.MMN2_g
+ N_XI1.XI7.NET27_XI1.XI7.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI7.MMN3 N_XI1.XI7.NET16_XI1.XI7.MMN3_d N_F_2_XI1.XI7.MMN3_g
+ N_XI1.XI7.NET28_XI1.XI7.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI7.MMinv2 N_BL<7>_XI1.XI7.MMinv2_d N_XI1.XI7.NET16_XI1.XI7.MMinv2_g
+ N_GND_XI1.XI7.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI7.MMinv2@4 N_BL<7>_XI1.XI7.MMinv2@4_d N_XI1.XI7.NET16_XI1.XI7.MMinv2@4_g
+ N_GND_XI1.XI7.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMinv2@3 N_BL<7>_XI1.XI7.MMinv2@3_d N_XI1.XI7.NET16_XI1.XI7.MMinv2@3_g
+ N_GND_XI1.XI7.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMinv2@2 N_BL<7>_XI1.XI7.MMinv2@2_d N_XI1.XI7.NET16_XI1.XI7.MMinv2@2_g
+ N_GND_XI1.XI7.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI7.MMP1 N_XI1.XI7.NET16_XI1.XI7.MMP1_d N_F_8_XI1.XI7.MMP1_g
+ N_VDD_XI1.XI7.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI7.MMP2 N_XI1.XI7.NET16_XI1.XI7.MMP2_d N_F_4_XI1.XI7.MMP2_g
+ N_VDD_XI1.XI7.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMP3 N_XI1.XI7.NET16_XI1.XI7.MMP3_d N_F_2_XI1.XI7.MMP3_g
+ N_VDD_XI1.XI7.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI7.MMen N_XI1.XI7.NET16_XI1.XI7.MMen_d N_EN_XI1.XI7.MMen_g
+ N_VDD_XI1.XI7.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI7.MMinv1 N_BL<7>_XI1.XI7.MMinv1_d N_XI1.XI7.NET16_XI1.XI7.MMinv1_g
+ N_VDD_XI1.XI7.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMinv1@4 N_BL<7>_XI1.XI7.MMinv1@4_d N_XI1.XI7.NET16_XI1.XI7.MMinv1@4_g
+ N_VDD_XI1.XI7.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMinv1@3 N_BL<7>_XI1.XI7.MMinv1@3_d N_XI1.XI7.NET16_XI1.XI7.MMinv1@3_g
+ N_VDD_XI1.XI7.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI7.MMinv1@2 N_BL<7>_XI1.XI7.MMinv1@2_d N_XI1.XI7.NET16_XI1.XI7.MMinv1@2_g
+ N_VDD_XI1.XI7.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI3.MMN1 N_XI1.XI3.NET27_XI1.XI3.MMN1_d N_F_8_INV_XI1.XI3.MMN1_g
+ N_GND_XI1.XI3.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI3.MMN2 N_XI1.XI3.NET28_XI1.XI3.MMN2_d N_F_4_XI1.XI3.MMN2_g
+ N_XI1.XI3.NET27_XI1.XI3.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI3.MMN3 N_XI1.XI3.NET16_XI1.XI3.MMN3_d N_F_2_XI1.XI3.MMN3_g
+ N_XI1.XI3.NET28_XI1.XI3.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI3.MMinv2 N_BL<3>_XI1.XI3.MMinv2_d N_XI1.XI3.NET16_XI1.XI3.MMinv2_g
+ N_GND_XI1.XI3.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI3.MMinv2@4 N_BL<3>_XI1.XI3.MMinv2@4_d N_XI1.XI3.NET16_XI1.XI3.MMinv2@4_g
+ N_GND_XI1.XI3.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMinv2@3 N_BL<3>_XI1.XI3.MMinv2@3_d N_XI1.XI3.NET16_XI1.XI3.MMinv2@3_g
+ N_GND_XI1.XI3.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMinv2@2 N_BL<3>_XI1.XI3.MMinv2@2_d N_XI1.XI3.NET16_XI1.XI3.MMinv2@2_g
+ N_GND_XI1.XI3.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI3.MMP1 N_XI1.XI3.NET16_XI1.XI3.MMP1_d N_F_8_INV_XI1.XI3.MMP1_g
+ N_VDD_XI1.XI3.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI3.MMP2 N_XI1.XI3.NET16_XI1.XI3.MMP2_d N_F_4_XI1.XI3.MMP2_g
+ N_VDD_XI1.XI3.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMP3 N_XI1.XI3.NET16_XI1.XI3.MMP3_d N_F_2_XI1.XI3.MMP3_g
+ N_VDD_XI1.XI3.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI3.MMen N_XI1.XI3.NET16_XI1.XI3.MMen_d N_EN_XI1.XI3.MMen_g
+ N_VDD_XI1.XI3.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI3.MMinv1 N_BL<3>_XI1.XI3.MMinv1_d N_XI1.XI3.NET16_XI1.XI3.MMinv1_g
+ N_VDD_XI1.XI3.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMinv1@4 N_BL<3>_XI1.XI3.MMinv1@4_d N_XI1.XI3.NET16_XI1.XI3.MMinv1@4_g
+ N_VDD_XI1.XI3.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMinv1@3 N_BL<3>_XI1.XI3.MMinv1@3_d N_XI1.XI3.NET16_XI1.XI3.MMinv1@3_g
+ N_VDD_XI1.XI3.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI3.MMinv1@2 N_BL<3>_XI1.XI3.MMinv1@2_d N_XI1.XI3.NET16_XI1.XI3.MMinv1@2_g
+ N_VDD_XI1.XI3.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI4.MMN1 N_XI1.XI4.NET27_XI1.XI4.MMN1_d N_F_8_XI1.XI4.MMN1_g
+ N_GND_XI1.XI4.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI4.MMN2 N_XI1.XI4.NET28_XI1.XI4.MMN2_d N_F_4_INV_XI1.XI4.MMN2_g
+ N_XI1.XI4.NET27_XI1.XI4.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI4.MMN3 N_XI1.XI4.NET16_XI1.XI4.MMN3_d N_F_2_INV_XI1.XI4.MMN3_g
+ N_XI1.XI4.NET28_XI1.XI4.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI4.MMinv2 N_BL<4>_XI1.XI4.MMinv2_d N_XI1.XI4.NET16_XI1.XI4.MMinv2_g
+ N_GND_XI1.XI4.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI4.MMinv2@4 N_BL<4>_XI1.XI4.MMinv2@4_d N_XI1.XI4.NET16_XI1.XI4.MMinv2@4_g
+ N_GND_XI1.XI4.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMinv2@3 N_BL<4>_XI1.XI4.MMinv2@3_d N_XI1.XI4.NET16_XI1.XI4.MMinv2@3_g
+ N_GND_XI1.XI4.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMinv2@2 N_BL<4>_XI1.XI4.MMinv2@2_d N_XI1.XI4.NET16_XI1.XI4.MMinv2@2_g
+ N_GND_XI1.XI4.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI4.MMP1 N_XI1.XI4.NET16_XI1.XI4.MMP1_d N_F_8_XI1.XI4.MMP1_g
+ N_VDD_XI1.XI4.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI4.MMP2 N_XI1.XI4.NET16_XI1.XI4.MMP2_d N_F_4_INV_XI1.XI4.MMP2_g
+ N_VDD_XI1.XI4.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMP3 N_XI1.XI4.NET16_XI1.XI4.MMP3_d N_F_2_INV_XI1.XI4.MMP3_g
+ N_VDD_XI1.XI4.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI4.MMen N_XI1.XI4.NET16_XI1.XI4.MMen_d N_EN_XI1.XI4.MMen_g
+ N_VDD_XI1.XI4.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI4.MMinv1 N_BL<4>_XI1.XI4.MMinv1_d N_XI1.XI4.NET16_XI1.XI4.MMinv1_g
+ N_VDD_XI1.XI4.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMinv1@4 N_BL<4>_XI1.XI4.MMinv1@4_d N_XI1.XI4.NET16_XI1.XI4.MMinv1@4_g
+ N_VDD_XI1.XI4.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMinv1@3 N_BL<4>_XI1.XI4.MMinv1@3_d N_XI1.XI4.NET16_XI1.XI4.MMinv1@3_g
+ N_VDD_XI1.XI4.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI4.MMinv1@2 N_BL<4>_XI1.XI4.MMinv1@2_d N_XI1.XI4.NET16_XI1.XI4.MMinv1@2_g
+ N_VDD_XI1.XI4.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI0.MMN1 N_XI1.XI0.NET27_XI1.XI0.MMN1_d N_F_8_INV_XI1.XI0.MMN1_g
+ N_GND_XI1.XI0.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI0.MMN2 N_XI1.XI0.NET28_XI1.XI0.MMN2_d N_F_4_INV_XI1.XI0.MMN2_g
+ N_XI1.XI0.NET27_XI1.XI0.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI0.MMN3 N_XI1.XI0.NET16_XI1.XI0.MMN3_d N_F_2_INV_XI1.XI0.MMN3_g
+ N_XI1.XI0.NET28_XI1.XI0.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI0.MMinv2 N_BL<0>_XI1.XI0.MMinv2_d N_XI1.XI0.NET16_XI1.XI0.MMinv2_g
+ N_GND_XI1.XI0.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI0.MMinv2@4 N_BL<0>_XI1.XI0.MMinv2@4_d N_XI1.XI0.NET16_XI1.XI0.MMinv2@4_g
+ N_GND_XI1.XI0.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMinv2@3 N_BL<0>_XI1.XI0.MMinv2@3_d N_XI1.XI0.NET16_XI1.XI0.MMinv2@3_g
+ N_GND_XI1.XI0.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMinv2@2 N_BL<0>_XI1.XI0.MMinv2@2_d N_XI1.XI0.NET16_XI1.XI0.MMinv2@2_g
+ N_GND_XI1.XI0.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI0.MMP1 N_XI1.XI0.NET16_XI1.XI0.MMP1_d N_F_8_INV_XI1.XI0.MMP1_g
+ N_VDD_XI1.XI0.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI0.MMP2 N_XI1.XI0.NET16_XI1.XI0.MMP2_d N_F_4_INV_XI1.XI0.MMP2_g
+ N_VDD_XI1.XI0.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMP3 N_XI1.XI0.NET16_XI1.XI0.MMP3_d N_F_2_INV_XI1.XI0.MMP3_g
+ N_VDD_XI1.XI0.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI0.MMen N_XI1.XI0.NET16_XI1.XI0.MMen_d N_EN_XI1.XI0.MMen_g
+ N_VDD_XI1.XI0.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI0.MMinv1 N_BL<0>_XI1.XI0.MMinv1_d N_XI1.XI0.NET16_XI1.XI0.MMinv1_g
+ N_VDD_XI1.XI0.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMinv1@4 N_BL<0>_XI1.XI0.MMinv1@4_d N_XI1.XI0.NET16_XI1.XI0.MMinv1@4_g
+ N_VDD_XI1.XI0.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMinv1@3 N_BL<0>_XI1.XI0.MMinv1@3_d N_XI1.XI0.NET16_XI1.XI0.MMinv1@3_g
+ N_VDD_XI1.XI0.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI0.MMinv1@2 N_BL<0>_XI1.XI0.MMinv1@2_d N_XI1.XI0.NET16_XI1.XI0.MMinv1@2_g
+ N_VDD_XI1.XI0.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI6.MMN1 N_XI1.XI6.NET27_XI1.XI6.MMN1_d N_F_8_XI1.XI6.MMN1_g
+ N_GND_XI1.XI6.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI6.MMN2 N_XI1.XI6.NET28_XI1.XI6.MMN2_d N_F_4_XI1.XI6.MMN2_g
+ N_XI1.XI6.NET27_XI1.XI6.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI6.MMN3 N_XI1.XI6.NET16_XI1.XI6.MMN3_d N_F_2_INV_XI1.XI6.MMN3_g
+ N_XI1.XI6.NET28_XI1.XI6.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI6.MMinv2 N_BL<6>_XI1.XI6.MMinv2_d N_XI1.XI6.NET16_XI1.XI6.MMinv2_g
+ N_GND_XI1.XI6.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI6.MMinv2@4 N_BL<6>_XI1.XI6.MMinv2@4_d N_XI1.XI6.NET16_XI1.XI6.MMinv2@4_g
+ N_GND_XI1.XI6.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMinv2@3 N_BL<6>_XI1.XI6.MMinv2@3_d N_XI1.XI6.NET16_XI1.XI6.MMinv2@3_g
+ N_GND_XI1.XI6.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMinv2@2 N_BL<6>_XI1.XI6.MMinv2@2_d N_XI1.XI6.NET16_XI1.XI6.MMinv2@2_g
+ N_GND_XI1.XI6.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI6.MMP1 N_XI1.XI6.NET16_XI1.XI6.MMP1_d N_F_8_XI1.XI6.MMP1_g
+ N_VDD_XI1.XI6.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI6.MMP2 N_XI1.XI6.NET16_XI1.XI6.MMP2_d N_F_4_XI1.XI6.MMP2_g
+ N_VDD_XI1.XI6.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMP3 N_XI1.XI6.NET16_XI1.XI6.MMP3_d N_F_2_INV_XI1.XI6.MMP3_g
+ N_VDD_XI1.XI6.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI6.MMen N_XI1.XI6.NET16_XI1.XI6.MMen_d N_EN_XI1.XI6.MMen_g
+ N_VDD_XI1.XI6.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI6.MMinv1 N_BL<6>_XI1.XI6.MMinv1_d N_XI1.XI6.NET16_XI1.XI6.MMinv1_g
+ N_VDD_XI1.XI6.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMinv1@4 N_BL<6>_XI1.XI6.MMinv1@4_d N_XI1.XI6.NET16_XI1.XI6.MMinv1@4_g
+ N_VDD_XI1.XI6.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMinv1@3 N_BL<6>_XI1.XI6.MMinv1@3_d N_XI1.XI6.NET16_XI1.XI6.MMinv1@3_g
+ N_VDD_XI1.XI6.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI6.MMinv1@2 N_BL<6>_XI1.XI6.MMinv1@2_d N_XI1.XI6.NET16_XI1.XI6.MMinv1@2_g
+ N_VDD_XI1.XI6.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI1.XI2.MMN1 N_XI1.XI2.NET27_XI1.XI2.MMN1_d N_F_8_INV_XI1.XI2.MMN1_g
+ N_GND_XI1.XI2.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=2.303e-13 PD=4.45e-07 PS=1.45e-06
mXI1.XI2.MMN2 N_XI1.XI2.NET28_XI1.XI2.MMN2_d N_F_4_XI1.XI2.MMN2_g
+ N_XI1.XI2.NET27_XI1.XI2.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.04575e-13 AS=1.04575e-13 PD=4.45e-07 PS=4.45e-07
mXI1.XI2.MMN3 N_XI1.XI2.NET16_XI1.XI2.MMN3_d N_F_2_INV_XI1.XI2.MMN3_g
+ N_XI1.XI2.NET28_XI1.XI2.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.538e-13 AS=1.04575e-13 PD=1.55e-06 PS=4.45e-07
mXI1.XI2.MMinv2 N_BL<2>_XI1.XI2.MMinv2_d N_XI1.XI2.NET16_XI1.XI2.MMinv2_g
+ N_GND_XI1.XI2.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07 AD=2.04e-13
+ AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI2.MMinv2@4 N_BL<2>_XI1.XI2.MMinv2@4_d N_XI1.XI2.NET16_XI1.XI2.MMinv2@4_g
+ N_GND_XI1.XI2.MMinv2@4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMinv2@3 N_BL<2>_XI1.XI2.MMinv2@3_d N_XI1.XI2.NET16_XI1.XI2.MMinv2@3_g
+ N_GND_XI1.XI2.MMinv2@3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=2.04e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMinv2@2 N_BL<2>_XI1.XI2.MMinv2@2_d N_XI1.XI2.NET16_XI1.XI2.MMinv2@2_g
+ N_GND_XI1.XI2.MMinv2@2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=8e-07
+ AD=2.04e-13 AS=3.92e-13 PD=5.1e-07 PS=1.78e-06
mXI1.XI2.MMP1 N_XI1.XI2.NET16_XI1.XI2.MMP1_d N_F_8_INV_XI1.XI2.MMP1_g
+ N_VDD_XI1.XI2.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=4.9e-13 PD=5.1e-07 PS=1.98e-06
mXI1.XI2.MMP2 N_XI1.XI2.NET16_XI1.XI2.MMP2_d N_F_4_XI1.XI2.MMP2_g
+ N_VDD_XI1.XI2.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06 AD=2.55e-13
+ AS=2.55e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMP3 N_XI1.XI2.NET16_XI1.XI2.MMP3_d N_F_2_INV_XI1.XI2.MMP3_g
+ N_VDD_XI1.XI2.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1e-06
+ AD=2.59091e-13 AS=2.55e-13 PD=5.54545e-07 PS=5.1e-07
mXI1.XI2.MMen N_XI1.XI2.NET16_XI1.XI2.MMen_d N_EN_XI1.XI2.MMen_g
+ N_VDD_XI1.XI2.MMen_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.10909e-13 AS=3.06e-13 PD=6.65455e-07 PS=5.1e-07
mXI1.XI2.MMinv1 N_BL<2>_XI1.XI2.MMinv1_d N_XI1.XI2.NET16_XI1.XI2.MMinv1_g
+ N_VDD_XI1.XI2.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMinv1@4 N_BL<2>_XI1.XI2.MMinv1@4_d N_XI1.XI2.NET16_XI1.XI2.MMinv1@4_g
+ N_VDD_XI1.XI2.MMinv1@4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMinv1@3 N_BL<2>_XI1.XI2.MMinv1@3_d N_XI1.XI2.NET16_XI1.XI2.MMinv1@3_g
+ N_VDD_XI1.XI2.MMinv1@3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=3.06e-13 PD=5.1e-07 PS=5.1e-07
mXI1.XI2.MMinv1@2 N_BL<2>_XI1.XI2.MMinv1@2_d N_XI1.XI2.NET16_XI1.XI2.MMinv1@2_g
+ N_VDD_XI1.XI2.MMinv1@2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=3.06e-13 AS=5.88e-13 PD=5.1e-07 PS=2.18e-06
mXI0.XI13.MMN1 N_XI0.XI13.NET14_XI0.XI13.MMN1_d N_F_32_XI0.XI13.MMN1_g
+ N_GND_XI0.XI13.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI14.MMN1 N_XI0.NET26_XI0.XI14.MMN1_d N_F_2_INV_XI0.XI14.MMN1_g
+ N_GND_XI0.XI14.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI13.MMN2 N_XI0.XI13.NET15_XI0.XI13.MMN2_d N_F_16_XI0.XI13.MMN2_g
+ N_XI0.XI13.NET14_XI0.XI13.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI14.MMN2 N_XI0.NET26_XI0.XI14.MMN2_d N_F_4_INV_XI0.XI14.MMN2_g
+ N_GND_XI0.XI14.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI13.MMN3 N_XI0.NET41_XI0.XI13.MMN3_d N_XI0.NET26_XI0.XI13.MMN3_g
+ N_XI0.XI13.NET15_XI0.XI13.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI14.MMN3 N_XI0.NET26_XI0.XI14.MMN3_d N_F_8_INV_XI0.XI14.MMN3_g
+ N_GND_XI0.XI14.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI13.MMP1 N_XI0.NET41_XI0.XI13.MMP1_d N_F_32_XI0.XI13.MMP1_g
+ N_VDD_XI0.XI13.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI14.MMP1 N_XI0.XI14.NET23_XI0.XI14.MMP1_d N_F_2_INV_XI0.XI14.MMP1_g
+ N_VDD_XI0.XI14.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI13.MMP2 N_XI0.NET41_XI0.XI13.MMP2_d N_F_16_XI0.XI13.MMP2_g
+ N_VDD_XI0.XI13.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI14.MMP2 N_XI0.XI14.NET24_XI0.XI14.MMP2_d N_F_4_INV_XI0.XI14.MMP2_g
+ N_XI0.XI14.NET23_XI0.XI14.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=2.4225e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI13.MMP3 N_XI0.NET41_XI0.XI13.MMP3_d N_XI0.NET26_XI0.XI13.MMP3_g
+ N_VDD_XI0.XI13.MMP3_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI14.MMP3 N_XI0.NET26_XI0.XI14.MMP3_d N_F_8_INV_XI0.XI14.MMP3_g
+ N_XI0.XI14.NET24_XI0.XI14.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI7.MMinv2 N_XI0.XI7.NET15_XI0.XI7.MMinv2_d N_XI0.NET32_XI0.XI7.MMinv2_g
+ N_GND_XI0.XI7.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI7.MMN3 N_X8.X12.noxref_9_XI0.XI7.MMN3_d N_XI0.NET32_XI0.XI7.MMN3_g
+ N_GND_XI0.XI7.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI7.MMN4 N_XI0.NET31_XI0.XI7.MMN4_d N_F_8_INV_XI0.XI7.MMN4_g
+ N_X8.X12.noxref_9_XI0.XI7.MMN4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI7.MMN2 N_XI0.NET31_XI0.XI7.MMN2_d N_XI0.XI7.NET15_XI0.XI7.MMN2_g
+ N_X8.X12.noxref_10_XI0.XI7.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI7.MMN1 N_X8.X12.noxref_10_XI0.XI7.MMN1_d N_F_8_XI0.XI7.MMN1_g
+ N_GND_XI0.XI7.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI7.MMinv1 N_XI0.XI7.NET15_XI0.XI7.MMinv1_d N_XI0.NET32_XI0.XI7.MMinv1_g
+ N_VDD_XI0.XI7.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI7.MMP3 N_X8.X12.noxref_8_XI0.XI7.MMP3_d N_XI0.NET32_XI0.XI7.MMP3_g
+ N_VDD_XI0.XI7.MMP3_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI7.MMP1 N_X8.X12.noxref_8_XI0.XI7.MMP1_d N_F_8_INV_XI0.XI7.MMP1_g
+ N_VDD_XI0.XI7.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI7.MMP4 N_XI0.NET31_XI0.XI7.MMP4_d N_XI0.XI7.NET15_XI0.XI7.MMP4_g
+ N_X8.X12.noxref_8_XI0.XI7.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI7.MMP2 N_XI0.NET31_XI0.XI7.MMP2_d N_F_8_XI0.XI7.MMP2_g
+ N_X8.X12.noxref_8_XI0.XI7.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI6.MMinv2 N_XI0.XI6.NET15_XI0.XI6.MMinv2_d N_F_2_XI0.XI6.MMinv2_g
+ N_GND_XI0.XI6.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI6.MMN3 N_X8.X13.noxref_9_XI0.XI6.MMN3_d N_F_2_XI0.XI6.MMN3_g
+ N_GND_XI0.XI6.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI6.MMN4 N_XI0.NET30_XI0.XI6.MMN4_d N_F_4_XI0.XI6.MMN4_g
+ N_X8.X13.noxref_9_XI0.XI6.MMN4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI6.MMN2 N_XI0.NET30_XI0.XI6.MMN2_d N_XI0.XI6.NET15_XI0.XI6.MMN2_g
+ N_X8.X13.noxref_10_XI0.XI6.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI6.MMN1 N_X8.X13.noxref_10_XI0.XI6.MMN1_d N_F_4_INV_XI0.XI6.MMN1_g
+ N_GND_XI0.XI6.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI6.MMinv1 N_XI0.XI6.NET15_XI0.XI6.MMinv1_d N_F_2_XI0.XI6.MMinv1_g
+ N_VDD_XI0.XI6.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI6.MMP3 N_X8.X13.noxref_8_XI0.XI6.MMP3_d N_F_2_XI0.XI6.MMP3_g
+ N_VDD_XI0.XI6.MMP3_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI6.MMP1 N_X8.X13.noxref_8_XI0.XI6.MMP1_d N_F_4_XI0.XI6.MMP1_g
+ N_VDD_XI0.XI6.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI6.MMP4 N_XI0.NET30_XI0.XI6.MMP4_d N_XI0.XI6.NET15_XI0.XI6.MMP4_g
+ N_X8.X13.noxref_8_XI0.XI6.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI6.MMP2 N_XI0.NET30_XI0.XI6.MMP2_d N_F_4_INV_XI0.XI6.MMP2_g
+ N_X8.X13.noxref_8_XI0.XI6.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI10.MMinv2 N_XI0.XI10.NET15_XI0.XI10.MMinv2_d
+ N_XI0.NET41_XI0.XI10.MMinv2_g N_GND_XI0.XI10.MMinv2_s N_GND_XI2.XI5.MMN1_b
+ N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI10.MMN3 N_X8.X14.noxref_9_XI0.XI10.MMN3_d N_XI0.NET41_XI0.XI10.MMN3_g
+ N_GND_XI0.XI10.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI10.MMN4 N_XI0.NET40_XI0.XI10.MMN4_d N_F_64_INV_XI0.XI10.MMN4_g
+ N_X8.X14.noxref_9_XI0.XI10.MMN4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI10.MMN2 N_XI0.NET40_XI0.XI10.MMN2_d N_XI0.XI10.NET15_XI0.XI10.MMN2_g
+ N_X8.X14.noxref_10_XI0.XI10.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI10.MMN1 N_X8.X14.noxref_10_XI0.XI10.MMN1_d N_F_64_XI0.XI10.MMN1_g
+ N_GND_XI0.XI10.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI10.MMinv1 N_XI0.XI10.NET15_XI0.XI10.MMinv1_d
+ N_XI0.NET41_XI0.XI10.MMinv1_g N_VDD_XI0.XI10.MMinv1_s N_VDD_XI0.XI7.MMinv1_b
+ P_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI10.MMP3 N_X8.X14.noxref_8_XI0.XI10.MMP3_d N_XI0.NET41_XI0.XI10.MMP3_g
+ N_VDD_XI0.XI10.MMP3_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI10.MMP1 N_X8.X14.noxref_8_XI0.XI10.MMP1_d N_F_64_INV_XI0.XI10.MMP1_g
+ N_VDD_XI0.XI10.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI10.MMP4 N_XI0.NET40_XI0.XI10.MMP4_d N_XI0.XI10.NET15_XI0.XI10.MMP4_g
+ N_X8.X14.noxref_8_XI0.XI10.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI10.MMP2 N_XI0.NET40_XI0.XI10.MMP2_d N_F_64_XI0.XI10.MMP2_g
+ N_X8.X14.noxref_8_XI0.XI10.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI9.MMinv2 N_XI0.XI9.NET15_XI0.XI9.MMinv2_d N_XI0.NET37_XI0.XI9.MMinv2_g
+ N_GND_XI0.XI9.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI9.MMN3 N_X8.X15.noxref_9_XI0.XI9.MMN3_d N_XI0.NET37_XI0.XI9.MMN3_g
+ N_GND_XI0.XI9.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI9.MMN4 N_XI0.NET36_XI0.XI9.MMN4_d N_F_32_INV_XI0.XI9.MMN4_g
+ N_X8.X15.noxref_9_XI0.XI9.MMN4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI9.MMN2 N_XI0.NET36_XI0.XI9.MMN2_d N_XI0.XI9.NET15_XI0.XI9.MMN2_g
+ N_X8.X15.noxref_10_XI0.XI9.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI9.MMN1 N_X8.X15.noxref_10_XI0.XI9.MMN1_d N_F_32_XI0.XI9.MMN1_g
+ N_GND_XI0.XI9.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI9.MMinv1 N_XI0.XI9.NET15_XI0.XI9.MMinv1_d N_XI0.NET37_XI0.XI9.MMinv1_g
+ N_VDD_XI0.XI9.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI9.MMP3 N_X8.X15.noxref_8_XI0.XI9.MMP3_d N_XI0.NET37_XI0.XI9.MMP3_g
+ N_VDD_XI0.XI9.MMP3_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI9.MMP1 N_X8.X15.noxref_8_XI0.XI9.MMP1_d N_F_32_INV_XI0.XI9.MMP1_g
+ N_VDD_XI0.XI9.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI9.MMP4 N_XI0.NET36_XI0.XI9.MMP4_d N_XI0.XI9.NET15_XI0.XI9.MMP4_g
+ N_X8.X15.noxref_8_XI0.XI9.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI9.MMP2 N_XI0.NET36_XI0.XI9.MMP2_d N_F_32_XI0.XI9.MMP2_g
+ N_X8.X15.noxref_8_XI0.XI9.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI8.MMinv2 N_XI0.XI8.NET15_XI0.XI8.MMinv2_d N_XI0.NET26_XI0.XI8.MMinv2_g
+ N_GND_XI0.XI8.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI8.MMN3 N_X8.X16.noxref_9_XI0.XI8.MMN3_d N_XI0.NET26_XI0.XI8.MMN3_g
+ N_GND_XI0.XI8.MMN3_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI8.MMN4 N_XI0.NET34_XI0.XI8.MMN4_d N_F_16_XI0.XI8.MMN4_g
+ N_X8.X16.noxref_9_XI0.XI8.MMN4_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI8.MMN2 N_XI0.NET34_XI0.XI8.MMN2_d N_XI0.XI8.NET15_XI0.XI8.MMN2_g
+ N_X8.X16.noxref_10_XI0.XI8.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07
+ W=4.7e-07 AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI8.MMN1 N_X8.X16.noxref_10_XI0.XI8.MMN1_d N_F_16_INV_XI0.XI8.MMN1_g
+ N_GND_XI0.XI8.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI8.MMinv1 N_XI0.XI8.NET15_XI0.XI8.MMinv1_d N_XI0.NET26_XI0.XI8.MMinv1_g
+ N_VDD_XI0.XI8.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI8.MMP3 N_X8.X16.noxref_8_XI0.XI8.MMP3_d N_XI0.NET26_XI0.XI8.MMP3_g
+ N_VDD_XI0.XI8.MMP3_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI8.MMP1 N_X8.X16.noxref_8_XI0.XI8.MMP1_d N_F_16_XI0.XI8.MMP1_g
+ N_VDD_XI0.XI8.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI8.MMP4 N_XI0.NET34_XI0.XI8.MMP4_d N_XI0.XI8.NET15_XI0.XI8.MMP4_g
+ N_X8.X16.noxref_8_XI0.XI8.MMP4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=1.1985e-13 PD=5.1e-07 PS=5.1e-07
mXI0.XI8.MMP2 N_XI0.NET34_XI0.XI8.MMP2_d N_F_16_INV_XI0.XI8.MMP2_g
+ N_X8.X16.noxref_8_XI0.XI8.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI11.MMN1 N_XI0.XI11.NET12_XI0.XI11.MMN1_d N_F_4_XI0.XI11.MMN1_g
+ N_GND_XI0.XI11.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI11.MMN2 N_XI0.NET32_XI0.XI11.MMN2_d N_F_2_XI0.XI11.MMN2_g
+ N_XI0.XI11.NET12_XI0.XI11.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI11.MMP1 N_XI0.NET32_XI0.XI11.MMP1_d N_F_4_XI0.XI11.MMP1_g
+ N_VDD_XI0.XI11.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI11.MMP2 N_XI0.NET32_XI0.XI11.MMP2_d N_F_2_XI0.XI11.MMP2_g
+ N_VDD_XI0.XI11.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI12.MMN1 N_XI0.XI12.NET12_XI0.XI12.MMN1_d N_F_16_XI0.XI12.MMN1_g
+ N_GND_XI0.XI12.MMN1_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI12.MMN2 N_XI0.NET37_XI0.XI12.MMN2_d N_XI0.NET26_XI0.XI12.MMN2_g
+ N_XI0.XI12.NET12_XI0.XI12.MMN2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI12.MMP1 N_XI0.NET37_XI0.XI12.MMP1_d N_F_16_XI0.XI12.MMP1_g
+ N_VDD_XI0.XI12.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI12.MMP2 N_XI0.NET37_XI0.XI12.MMP2_d N_XI0.NET26_XI0.XI12.MMP2_g
+ N_VDD_XI0.XI12.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI2.MM0 N_XI0.XI2.NET16_XI0.XI2.MM0_d N_XI0.NET31_XI0.XI2.MM0_g
+ N_GND_XI0.XI2.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI2.MMN5 N_XI0.XI2.NET20_XI0.XI2.MMN5_d N_XI0.XI2.NET16_XI0.XI2.MMN5_g
+ N_XI0.XI2.NET37_XI0.XI2.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI2.MMN6 N_XI0.XI2.NET37_XI0.XI2.MMN6_d N_CLK_IN_XI0.XI2.MMN6_g
+ N_GND_XI0.XI2.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI2.MMN8 N_F_8_INV_XI0.XI2.MMN8_d N_CLK_IN_XI0.XI2.MMN8_g
+ N_XI0.XI2.NET36_XI0.XI2.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI2.MMN9 N_XI0.XI2.NET36_XI0.XI2.MMN9_d N_XI0.XI2.NET20_XI0.XI2.MMN9_g
+ N_GND_XI0.XI2.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI2.MMinv2 N_F_8_XI0.XI2.MMinv2_d N_F_8_INV_XI0.XI2.MMinv2_g
+ N_GND_XI0.XI2.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI2.MMP1 N_XI0.XI2.NET38_XI0.XI2.MMP1_d N_XI0.NET31_XI0.XI2.MMP1_g
+ N_VDD_XI0.XI2.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI2.MMP2 N_XI0.XI2.NET16_XI0.XI2.MMP2_d N_CLK_IN_XI0.XI2.MMP2_g
+ N_XI0.XI2.NET38_XI0.XI2.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI2.MMP4 N_XI0.XI2.NET20_XI0.XI2.MMP4_d N_CLK_IN_XI0.XI2.MMP4_g
+ N_VDD_XI0.XI2.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI2.MMP7 N_F_8_INV_XI0.XI2.MMP7_d N_XI0.XI2.NET20_XI0.XI2.MMP7_g
+ N_VDD_XI0.XI2.MMP7_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI2.MMrst N_F_8_INV_XI0.XI2.MMrst_d N_RST_XI0.XI2.MMrst_g
+ N_VDD_XI0.XI2.MMrst_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI2.MMinv1 N_F_8_XI0.XI2.MMinv1_d N_F_8_INV_XI0.XI2.MMinv1_g
+ N_VDD_XI0.XI2.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI1.MM0 N_XI0.XI1.NET16_XI0.XI1.MM0_d N_XI0.NET30_XI0.XI1.MM0_g
+ N_GND_XI0.XI1.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI1.MMN5 N_XI0.XI1.NET20_XI0.XI1.MMN5_d N_XI0.XI1.NET16_XI0.XI1.MMN5_g
+ N_XI0.XI1.NET37_XI0.XI1.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI1.MMN6 N_XI0.XI1.NET37_XI0.XI1.MMN6_d N_CLK_IN_XI0.XI1.MMN6_g
+ N_GND_XI0.XI1.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI1.MMN8 N_F_4_INV_XI0.XI1.MMN8_d N_CLK_IN_XI0.XI1.MMN8_g
+ N_XI0.XI1.NET36_XI0.XI1.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI1.MMN9 N_XI0.XI1.NET36_XI0.XI1.MMN9_d N_XI0.XI1.NET20_XI0.XI1.MMN9_g
+ N_GND_XI0.XI1.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI1.MMinv2 N_F_4_XI0.XI1.MMinv2_d N_F_4_INV_XI0.XI1.MMinv2_g
+ N_GND_XI0.XI1.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI1.MMP1 N_XI0.XI1.NET38_XI0.XI1.MMP1_d N_XI0.NET30_XI0.XI1.MMP1_g
+ N_VDD_XI0.XI1.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI1.MMP2 N_XI0.XI1.NET16_XI0.XI1.MMP2_d N_CLK_IN_XI0.XI1.MMP2_g
+ N_XI0.XI1.NET38_XI0.XI1.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI1.MMP4 N_XI0.XI1.NET20_XI0.XI1.MMP4_d N_CLK_IN_XI0.XI1.MMP4_g
+ N_VDD_XI0.XI1.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI1.MMP7 N_F_4_INV_XI0.XI1.MMP7_d N_XI0.XI1.NET20_XI0.XI1.MMP7_g
+ N_VDD_XI0.XI1.MMP7_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI1.MMrst N_F_4_INV_XI0.XI1.MMrst_d N_RST_XI0.XI1.MMrst_g
+ N_VDD_XI0.XI1.MMrst_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI1.MMinv1 N_F_4_XI0.XI1.MMinv1_d N_F_4_INV_XI0.XI1.MMinv1_g
+ N_VDD_XI0.XI1.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI0.MM0 N_XI0.XI0.NET16_XI0.XI0.MM0_d N_F_2_INV_XI0.XI0.MM0_g
+ N_GND_XI0.XI0.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI0.MMN5 N_XI0.XI0.NET20_XI0.XI0.MMN5_d N_XI0.XI0.NET16_XI0.XI0.MMN5_g
+ N_XI0.XI0.NET37_XI0.XI0.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI0.MMN6 N_XI0.XI0.NET37_XI0.XI0.MMN6_d N_CLK_IN_XI0.XI0.MMN6_g
+ N_GND_XI0.XI0.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI0.MMN8 N_F_2_INV_XI0.XI0.MMN8_d N_CLK_IN_XI0.XI0.MMN8_g
+ N_XI0.XI0.NET36_XI0.XI0.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI0.MMN9 N_XI0.XI0.NET36_XI0.XI0.MMN9_d N_XI0.XI0.NET20_XI0.XI0.MMN9_g
+ N_GND_XI0.XI0.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI0.MMinv2 N_F_2_XI0.XI0.MMinv2_d N_F_2_INV_XI0.XI0.MMinv2_g
+ N_GND_XI0.XI0.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI0.MMP1 N_XI0.XI0.NET38_XI0.XI0.MMP1_d N_F_2_INV_XI0.XI0.MMP1_g
+ N_VDD_XI0.XI0.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI0.MMP2 N_XI0.XI0.NET16_XI0.XI0.MMP2_d N_CLK_IN_XI0.XI0.MMP2_g
+ N_XI0.XI0.NET38_XI0.XI0.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI0.MMP4 N_XI0.XI0.NET20_XI0.XI0.MMP4_d N_CLK_IN_XI0.XI0.MMP4_g
+ N_VDD_XI0.XI0.MMP4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI0.MMP7 N_F_2_INV_XI0.XI0.MMP7_d N_XI0.XI0.NET20_XI0.XI0.MMP7_g
+ N_VDD_XI0.XI0.MMP7_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI0.MMrst N_F_2_INV_XI0.XI0.MMrst_d N_RST_XI0.XI0.MMrst_g
+ N_VDD_XI0.XI0.MMrst_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI0.MMinv1 N_F_2_XI0.XI0.MMinv1_d N_F_2_INV_XI0.XI0.MMinv1_g
+ N_VDD_XI0.XI0.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI5.MM0 N_XI0.XI5.NET16_XI0.XI5.MM0_d N_XI0.NET40_XI0.XI5.MM0_g
+ N_GND_XI0.XI5.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI5.MMN5 N_XI0.XI5.NET20_XI0.XI5.MMN5_d N_XI0.XI5.NET16_XI0.XI5.MMN5_g
+ N_XI0.XI5.NET37_XI0.XI5.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI5.MMN6 N_XI0.XI5.NET37_XI0.XI5.MMN6_d N_CLK_IN_XI0.XI5.MMN6_g
+ N_GND_XI0.XI5.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI5.MMN8 N_F_64_INV_XI0.XI5.MMN8_d N_CLK_IN_XI0.XI5.MMN8_g
+ N_XI0.XI5.NET36_XI0.XI5.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI5.MMN9 N_XI0.XI5.NET36_XI0.XI5.MMN9_d N_XI0.XI5.NET20_XI0.XI5.MMN9_g
+ N_GND_XI0.XI5.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI5.MMinv2 N_F_64_XI0.XI5.MMinv2_d N_F_64_INV_XI0.XI5.MMinv2_g
+ N_GND_XI0.XI5.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI5.MMP1 N_XI0.XI5.NET38_XI0.XI5.MMP1_d N_XI0.NET40_XI0.XI5.MMP1_g
+ N_VDD_XI0.XI5.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI5.MMP2 N_XI0.XI5.NET16_XI0.XI5.MMP2_d N_CLK_IN_XI0.XI5.MMP2_g
+ N_XI0.XI5.NET38_XI0.XI5.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI5.MMP4 N_XI0.XI5.NET20_XI0.XI5.MMP4_d N_CLK_IN_XI0.XI5.MMP4_g
+ N_VDD_XI0.XI5.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI5.MMP7 N_F_64_INV_XI0.XI5.MMP7_d N_XI0.XI5.NET20_XI0.XI5.MMP7_g
+ N_VDD_XI0.XI5.MMP7_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI5.MMrst N_F_64_INV_XI0.XI5.MMrst_d N_RST_XI0.XI5.MMrst_g
+ N_VDD_XI0.XI5.MMrst_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI5.MMinv1 N_F_64_XI0.XI5.MMinv1_d N_F_64_INV_XI0.XI5.MMinv1_g
+ N_VDD_XI0.XI5.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI4.MM0 N_XI0.XI4.NET16_XI0.XI4.MM0_d N_XI0.NET36_XI0.XI4.MM0_g
+ N_GND_XI0.XI4.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI4.MMN5 N_XI0.XI4.NET20_XI0.XI4.MMN5_d N_XI0.XI4.NET16_XI0.XI4.MMN5_g
+ N_XI0.XI4.NET37_XI0.XI4.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI4.MMN6 N_XI0.XI4.NET37_XI0.XI4.MMN6_d N_CLK_IN_XI0.XI4.MMN6_g
+ N_GND_XI0.XI4.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI4.MMN8 N_F_32_INV_XI0.XI4.MMN8_d N_CLK_IN_XI0.XI4.MMN8_g
+ N_XI0.XI4.NET36_XI0.XI4.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI4.MMN9 N_XI0.XI4.NET36_XI0.XI4.MMN9_d N_XI0.XI4.NET20_XI0.XI4.MMN9_g
+ N_GND_XI0.XI4.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI4.MMinv2 N_F_32_XI0.XI4.MMinv2_d N_F_32_INV_XI0.XI4.MMinv2_g
+ N_GND_XI0.XI4.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI4.MMP1 N_XI0.XI4.NET38_XI0.XI4.MMP1_d N_XI0.NET36_XI0.XI4.MMP1_g
+ N_VDD_XI0.XI4.MMP1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI4.MMP2 N_XI0.XI4.NET16_XI0.XI4.MMP2_d N_CLK_IN_XI0.XI4.MMP2_g
+ N_XI0.XI4.NET38_XI0.XI4.MMP2_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI4.MMP4 N_XI0.XI4.NET20_XI0.XI4.MMP4_d N_CLK_IN_XI0.XI4.MMP4_g
+ N_VDD_XI0.XI4.MMP4_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI4.MMP7 N_F_32_INV_XI0.XI4.MMP7_d N_XI0.XI4.NET20_XI0.XI4.MMP7_g
+ N_VDD_XI0.XI4.MMP7_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI4.MMrst N_F_32_INV_XI0.XI4.MMrst_d N_RST_XI0.XI4.MMrst_g
+ N_VDD_XI0.XI4.MMrst_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI4.MMinv1 N_F_32_XI0.XI4.MMinv1_d N_F_32_INV_XI0.XI4.MMinv1_g
+ N_VDD_XI0.XI4.MMinv1_s N_VDD_XI0.XI7.MMinv1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI3.MM0 N_XI0.XI3.NET16_XI0.XI3.MM0_d N_XI0.NET34_XI0.XI3.MM0_g
+ N_GND_XI0.XI3.MM0_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07 AD=2.303e-13
+ AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI3.MMN5 N_XI0.XI3.NET20_XI0.XI3.MMN5_d N_XI0.XI3.NET16_XI0.XI3.MMN5_g
+ N_XI0.XI3.NET37_XI0.XI3.MMN5_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI3.MMN6 N_XI0.XI3.NET37_XI0.XI3.MMN6_d N_CLK_IN_XI0.XI3.MMN6_g
+ N_GND_XI0.XI3.MMN6_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI3.MMN8 N_F_16_INV_XI0.XI3.MMN8_d N_CLK_IN_XI0.XI3.MMN8_g
+ N_XI0.XI3.NET36_XI0.XI3.MMN8_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=1.1985e-13 PD=1.45e-06 PS=5.1e-07
mXI0.XI3.MMN9 N_XI0.XI3.NET36_XI0.XI3.MMN9_d N_XI0.XI3.NET20_XI0.XI3.MMN9_g
+ N_GND_XI0.XI3.MMN9_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=1.1985e-13 AS=2.303e-13 PD=5.1e-07 PS=1.45e-06
mXI0.XI3.MMinv2 N_F_16_XI0.XI3.MMinv2_d N_F_16_INV_XI0.XI3.MMinv2_g
+ N_GND_XI0.XI3.MMinv2_s N_GND_XI2.XI5.MMN1_b N_18 L=1.8e-07 W=4.7e-07
+ AD=2.303e-13 AS=2.303e-13 PD=1.45e-06 PS=1.45e-06
mXI0.XI3.MMP1 N_XI0.XI3.NET38_XI0.XI3.MMP1_d N_XI0.NET34_XI0.XI3.MMP1_g
+ N_VDD_XI0.XI3.MMP1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=2.4225e-13 AS=4.655e-13 PD=5.1e-07 PS=1.93e-06
mXI0.XI3.MMP2 N_XI0.XI3.NET16_XI0.XI3.MMP2_d N_CLK_IN_XI0.XI3.MMP2_g
+ N_XI0.XI3.NET38_XI0.XI3.MMP2_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=2.4225e-13 PD=1.93e-06 PS=5.1e-07
mXI0.XI3.MMP4 N_XI0.XI3.NET20_XI0.XI3.MMP4_d N_CLK_IN_XI0.XI3.MMP4_g
+ N_VDD_XI0.XI3.MMP4_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI3.MMP7 N_F_16_INV_XI0.XI3.MMP7_d N_XI0.XI3.NET20_XI0.XI3.MMP7_g
+ N_VDD_XI0.XI3.MMP7_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
mXI0.XI3.MMrst N_F_16_INV_XI0.XI3.MMrst_d N_RST_XI0.XI3.MMrst_g
+ N_VDD_XI0.XI3.MMrst_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=1.2e-06
+ AD=5.88e-13 AS=5.88e-13 PD=2.18e-06 PS=2.18e-06
mXI0.XI3.MMinv1 N_F_16_XI0.XI3.MMinv1_d N_F_16_INV_XI0.XI3.MMinv1_g
+ N_VDD_XI0.XI3.MMinv1_s N_VDD_XI2.XI5.MMP1_b P_18 L=1.8e-07 W=9.5e-07
+ AD=4.655e-13 AS=4.655e-13 PD=1.93e-06 PS=1.93e-06
*
.include "total.pex.spi.TOTAL.pxi"
*
.ends
*
*
