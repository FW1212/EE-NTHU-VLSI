* File: clkgen.pex.spi
* Created: Mon Oct 30 21:28:24 2023
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "clkgen.pex.spi.pex"
.subckt clkgen  TRIGGER CLKOUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* CLKOUT	CLKOUT
* TRIGGER	TRIGGER
mXI1.MM0 N_NET15_XI1.MM0_d N_TRIGGER_XI1.MM0_g N_XI1.NET18_XI1.MM0_s
+ N_VSS_XI2.MM1_b N_18 L=2e-07 W=2e-06 AD=9.8e-13 AS=5.1e-13 PD=2.98e-06
+ PS=5.1e-07
mXI1.MM1 N_XI1.NET18_XI1.MM1_d N_CLKOUT_XI1.MM1_g N_VSS_XI1.MM1_s
+ N_VSS_XI2.MM1_b N_18 L=2e-07 W=2e-06 AD=5.1e-13 AS=9.8e-13 PD=5.1e-07
+ PS=2.98e-06
mXI1.MM2 N_NET15_XI1.MM2_d N_TRIGGER_XI1.MM2_g N_VDD_XI1.MM2_s N_VDD_XI2.MM0_b
+ P_18 L=2e-07 W=3e-06 AD=7.65e-13 AS=1.47e-12 PD=5.1e-07 PS=3.98e-06
mXI1.MM3 N_NET15_XI1.MM3_d N_CLKOUT_XI1.MM3_g N_VDD_XI1.MM3_s N_VDD_XI2.MM0_b
+ P_18 L=2e-07 W=3e-06 AD=7.65e-13 AS=1.47e-12 PD=5.1e-07 PS=3.98e-06
mXI2.MM1 N_NET14_XI2.MM1_d N_NET15_XI2.MM1_g N_VSS_XI2.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI2.MM0 N_NET14_XI2.MM0_d N_NET15_XI2.MM0_g N_VDD_XI2.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI3.MM1 N_NET13_XI3.MM1_d N_NET14_XI3.MM1_g N_VSS_XI3.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI3.MM0 N_NET13_XI3.MM0_d N_NET14_XI3.MM0_g N_VDD_XI3.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI4.MM1 N_NET12_XI4.MM1_d N_NET13_XI4.MM1_g N_VSS_XI4.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI4.MM0 N_NET12_XI4.MM0_d N_NET13_XI4.MM0_g N_VDD_XI4.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI5.MM1 N_NET11_XI5.MM1_d N_NET12_XI5.MM1_g N_VSS_XI5.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI5.MM0 N_NET11_XI5.MM0_d N_NET12_XI5.MM0_g N_VDD_XI5.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI6.MM1 N_NET10_XI6.MM1_d N_NET11_XI6.MM1_g N_VSS_XI6.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI6.MM0 N_NET10_XI6.MM0_d N_NET11_XI6.MM0_g N_VDD_XI6.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
mXI7.MM1 N_CLKOUT_XI7.MM1_d N_NET10_XI7.MM1_g N_VSS_XI7.MM1_s N_VSS_XI2.MM1_b
+ N_18 L=1.8e-07 W=1e-06 AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
mXI7.MM0 N_CLKOUT_XI7.MM0_d N_NET10_XI7.MM0_g N_VDD_XI7.MM0_s N_VDD_XI2.MM0_b
+ P_18 L=1.8e-07 W=3e-06 AD=1.47e-12 AS=1.47e-12 PD=3.98e-06 PS=3.98e-06
*
.include "clkgen.pex.spi.CLKGEN.pxi"
*
.ends
*
*
