* File: buf.pex.spi
* Created: Mon Oct 30 15:23:23 2023
* Program "Calibre xRC"
* Version "v2016.4_15.11"
* 
.include "buf.pex.spi.pex"
.subckt buf  A OUT VSS VDD
* 
* VDD	VDD
* VSS	VSS
* OUT	OUT
* A	A
MM2 N_NET12_MM2_d N_A_MM2_g N_VSS_MM2_s N_VSS_MM2_b N_18 L=1.8e-07 W=5e-07
+ AD=2.45e-13 AS=2.45e-13 PD=1.48e-06 PS=1.48e-06
MM4 N_OUT_MM4_d N_NET12_MM4_g N_VSS_MM4_s N_VSS_MM2_b N_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
MM1 N_NET12_MM1_d N_A_MM1_g N_VDD_MM1_s N_VDD_MM1_b P_18 L=1.8e-07 W=1e-06
+ AD=4.9e-13 AS=4.9e-13 PD=1.98e-06 PS=1.98e-06
MM3 N_OUT_MM3_d N_NET12_MM3_g N_VDD_MM3_s N_VDD_MM1_b P_18 L=1.8e-07 W=2.67e-06
+ AD=1.3083e-12 AS=1.3083e-12 PD=3.65e-06 PS=3.65e-06
*
.include "buf.pex.spi.BUF.pxi"
*
.ends
*
*
