************************************************************************
* auCdl Netlist:
* 
* Library Name:  323002mylib
* Top Cell Name: inv
* View Name:     schematic
* Netlisted on:  Sep 28 20:50:15 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: 323002mylib
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv A Out VDD VSS
*.PININFO A:I VDD:I VSS:I Out:O
MM0 Out A VDD VDD p_18 W=3u L=180.00n
MM1 Out A VSS VSS n_18 W=1u L=180.00n
.ENDS

