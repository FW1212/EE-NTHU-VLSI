************************************************************************
* auCdl Netlist:
* 
* Library Name:  323002mylib
* Top Cell Name: clkgen
* View Name:     schematic
* Netlisted on:  Oct  4 02:06:16 2023
************************************************************************

*.BIPOLAR
*.RESI = 2000 
*.RESVAL
*.CAPVAL
*.DIOPERI
*.DIOAREA
*.EQUATION
*.SCALE METER
*.MEGA
.PARAM



************************************************************************
* Library Name: 323002mylib
* Cell Name:    nand2
* View Name:    schematic
************************************************************************

.SUBCKT nand2 A B Vdd Vout Vss
*.PININFO A:I B:I Vdd:I Vss:I Vout:O
MM1 net18 B Vss Vss n_18 W=2u L=200.0n
MM0 Vout A net18 Vss n_18 W=2u L=200.0n
MM3 Vout B Vdd Vdd p_18 W=3u L=200.0n
MM2 Vout A Vdd Vdd p_18 W=3u L=200.0n
.ENDS

************************************************************************
* Library Name: 323002mylib
* Cell Name:    inv
* View Name:    schematic
************************************************************************

.SUBCKT inv A Out VDD VSS
*.PININFO A:I VDD:I VSS:I Out:O
MM0 Out A VDD VDD p_18 W=3u L=180.00n
MM1 Out A VSS VSS n_18 W=1u L=180.00n
.ENDS

************************************************************************
* Library Name: 323002mylib
* Cell Name:    clkgen
* View Name:    schematic
************************************************************************

.SUBCKT clkgen Vdd Vss clkout trigger
*.PININFO Vdd:I Vss:I trigger:I clkout:O
XNAND0 trigger clkout Vdd net15 Vss / nand2
Xinv5 net10 clkout Vdd Vss / inv
Xinv4 net11 net10 Vdd Vss / inv
Xinv3 net12 net11 Vdd Vss / inv
Xinv2 net13 net12 Vdd Vss / inv
Xinv1 net14 net13 Vdd Vss / inv
Xinv0 net15 net14 Vdd Vss / inv
.ENDS

